magic
tech sky130A
magscale 1 2
timestamp 1634569069
<< obsli1 >>
rect 1104 2159 59403 37553
<< obsm1 >>
rect 198 2128 59878 38616
<< metal2 >>
rect 202 39200 258 40000
rect 662 39200 718 40000
rect 1214 39200 1270 40000
rect 1766 39200 1822 40000
rect 2226 39200 2282 40000
rect 2778 39200 2834 40000
rect 3330 39200 3386 40000
rect 3882 39200 3938 40000
rect 4342 39200 4398 40000
rect 4894 39200 4950 40000
rect 5446 39200 5502 40000
rect 5906 39200 5962 40000
rect 6458 39200 6514 40000
rect 7010 39200 7066 40000
rect 7562 39200 7618 40000
rect 8022 39200 8078 40000
rect 8574 39200 8630 40000
rect 9126 39200 9182 40000
rect 9586 39200 9642 40000
rect 10138 39200 10194 40000
rect 10690 39200 10746 40000
rect 11242 39200 11298 40000
rect 11702 39200 11758 40000
rect 12254 39200 12310 40000
rect 12806 39200 12862 40000
rect 13266 39200 13322 40000
rect 13818 39200 13874 40000
rect 14370 39200 14426 40000
rect 14922 39200 14978 40000
rect 15382 39200 15438 40000
rect 15934 39200 15990 40000
rect 16486 39200 16542 40000
rect 17038 39200 17094 40000
rect 17498 39200 17554 40000
rect 18050 39200 18106 40000
rect 18602 39200 18658 40000
rect 19062 39200 19118 40000
rect 19614 39200 19670 40000
rect 20166 39200 20222 40000
rect 20718 39200 20774 40000
rect 21178 39200 21234 40000
rect 21730 39200 21786 40000
rect 22282 39200 22338 40000
rect 22742 39200 22798 40000
rect 23294 39200 23350 40000
rect 23846 39200 23902 40000
rect 24398 39200 24454 40000
rect 24858 39200 24914 40000
rect 25410 39200 25466 40000
rect 25962 39200 26018 40000
rect 26422 39200 26478 40000
rect 26974 39200 27030 40000
rect 27526 39200 27582 40000
rect 28078 39200 28134 40000
rect 28538 39200 28594 40000
rect 29090 39200 29146 40000
rect 29642 39200 29698 40000
rect 30194 39200 30250 40000
rect 30654 39200 30710 40000
rect 31206 39200 31262 40000
rect 31758 39200 31814 40000
rect 32218 39200 32274 40000
rect 32770 39200 32826 40000
rect 33322 39200 33378 40000
rect 33874 39200 33930 40000
rect 34334 39200 34390 40000
rect 34886 39200 34942 40000
rect 35438 39200 35494 40000
rect 35898 39200 35954 40000
rect 36450 39200 36506 40000
rect 37002 39200 37058 40000
rect 37554 39200 37610 40000
rect 38014 39200 38070 40000
rect 38566 39200 38622 40000
rect 39118 39200 39174 40000
rect 39578 39200 39634 40000
rect 40130 39200 40186 40000
rect 40682 39200 40738 40000
rect 41234 39200 41290 40000
rect 41694 39200 41750 40000
rect 42246 39200 42302 40000
rect 42798 39200 42854 40000
rect 43258 39200 43314 40000
rect 43810 39200 43866 40000
rect 44362 39200 44418 40000
rect 44914 39200 44970 40000
rect 45374 39200 45430 40000
rect 45926 39200 45982 40000
rect 46478 39200 46534 40000
rect 47030 39200 47086 40000
rect 47490 39200 47546 40000
rect 48042 39200 48098 40000
rect 48594 39200 48650 40000
rect 49054 39200 49110 40000
rect 49606 39200 49662 40000
rect 50158 39200 50214 40000
rect 50710 39200 50766 40000
rect 51170 39200 51226 40000
rect 51722 39200 51778 40000
rect 52274 39200 52330 40000
rect 52734 39200 52790 40000
rect 53286 39200 53342 40000
rect 53838 39200 53894 40000
rect 54390 39200 54446 40000
rect 54850 39200 54906 40000
rect 55402 39200 55458 40000
rect 55954 39200 56010 40000
rect 56414 39200 56470 40000
rect 56966 39200 57022 40000
rect 57518 39200 57574 40000
rect 58070 39200 58126 40000
rect 58530 39200 58586 40000
rect 59082 39200 59138 40000
rect 59634 39200 59690 40000
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 294 0 350 800
rect 478 0 534 800
rect 570 0 626 800
rect 662 0 718 800
rect 846 0 902 800
rect 938 0 994 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57886 0 57942 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 58990 0 59046 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59358 0 59414 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59726 0 59782 800
rect 59818 0 59874 800
<< obsm2 >>
rect 314 39144 606 39250
rect 774 39144 1158 39250
rect 1326 39144 1710 39250
rect 1878 39144 2170 39250
rect 2338 39144 2722 39250
rect 2890 39144 3274 39250
rect 3442 39144 3826 39250
rect 3994 39144 4286 39250
rect 4454 39144 4838 39250
rect 5006 39144 5390 39250
rect 5558 39144 5850 39250
rect 6018 39144 6402 39250
rect 6570 39144 6954 39250
rect 7122 39144 7506 39250
rect 7674 39144 7966 39250
rect 8134 39144 8518 39250
rect 8686 39144 9070 39250
rect 9238 39144 9530 39250
rect 9698 39144 10082 39250
rect 10250 39144 10634 39250
rect 10802 39144 11186 39250
rect 11354 39144 11646 39250
rect 11814 39144 12198 39250
rect 12366 39144 12750 39250
rect 12918 39144 13210 39250
rect 13378 39144 13762 39250
rect 13930 39144 14314 39250
rect 14482 39144 14866 39250
rect 15034 39144 15326 39250
rect 15494 39144 15878 39250
rect 16046 39144 16430 39250
rect 16598 39144 16982 39250
rect 17150 39144 17442 39250
rect 17610 39144 17994 39250
rect 18162 39144 18546 39250
rect 18714 39144 19006 39250
rect 19174 39144 19558 39250
rect 19726 39144 20110 39250
rect 20278 39144 20662 39250
rect 20830 39144 21122 39250
rect 21290 39144 21674 39250
rect 21842 39144 22226 39250
rect 22394 39144 22686 39250
rect 22854 39144 23238 39250
rect 23406 39144 23790 39250
rect 23958 39144 24342 39250
rect 24510 39144 24802 39250
rect 24970 39144 25354 39250
rect 25522 39144 25906 39250
rect 26074 39144 26366 39250
rect 26534 39144 26918 39250
rect 27086 39144 27470 39250
rect 27638 39144 28022 39250
rect 28190 39144 28482 39250
rect 28650 39144 29034 39250
rect 29202 39144 29586 39250
rect 29754 39144 30138 39250
rect 30306 39144 30598 39250
rect 30766 39144 31150 39250
rect 31318 39144 31702 39250
rect 31870 39144 32162 39250
rect 32330 39144 32714 39250
rect 32882 39144 33266 39250
rect 33434 39144 33818 39250
rect 33986 39144 34278 39250
rect 34446 39144 34830 39250
rect 34998 39144 35382 39250
rect 35550 39144 35842 39250
rect 36010 39144 36394 39250
rect 36562 39144 36946 39250
rect 37114 39144 37498 39250
rect 37666 39144 37958 39250
rect 38126 39144 38510 39250
rect 38678 39144 39062 39250
rect 39230 39144 39522 39250
rect 39690 39144 40074 39250
rect 40242 39144 40626 39250
rect 40794 39144 41178 39250
rect 41346 39144 41638 39250
rect 41806 39144 42190 39250
rect 42358 39144 42742 39250
rect 42910 39144 43202 39250
rect 43370 39144 43754 39250
rect 43922 39144 44306 39250
rect 44474 39144 44858 39250
rect 45026 39144 45318 39250
rect 45486 39144 45870 39250
rect 46038 39144 46422 39250
rect 46590 39144 46974 39250
rect 47142 39144 47434 39250
rect 47602 39144 47986 39250
rect 48154 39144 48538 39250
rect 48706 39144 48998 39250
rect 49166 39144 49550 39250
rect 49718 39144 50102 39250
rect 50270 39144 50654 39250
rect 50822 39144 51114 39250
rect 51282 39144 51666 39250
rect 51834 39144 52218 39250
rect 52386 39144 52678 39250
rect 52846 39144 53230 39250
rect 53398 39144 53782 39250
rect 53950 39144 54334 39250
rect 54502 39144 54794 39250
rect 54962 39144 55346 39250
rect 55514 39144 55898 39250
rect 56066 39144 56358 39250
rect 56526 39144 56910 39250
rect 57078 39144 57462 39250
rect 57630 39144 58014 39250
rect 58182 39144 58474 39250
rect 58642 39144 59026 39250
rect 59194 39144 59578 39250
rect 59746 39144 59872 39250
rect 204 856 59872 39144
rect 406 800 422 856
rect 774 800 790 856
rect 1142 800 1158 856
rect 1510 800 1526 856
rect 1878 800 1894 856
rect 2246 800 2262 856
rect 2614 800 2630 856
rect 2982 800 2998 856
rect 3350 800 3366 856
rect 3810 800 3826 856
rect 4178 800 4194 856
rect 4546 800 4562 856
rect 4914 800 4930 856
rect 5282 800 5298 856
rect 5650 800 5666 856
rect 6018 800 6034 856
rect 6386 800 6402 856
rect 6754 800 6770 856
rect 7122 800 7138 856
rect 7582 800 7598 856
rect 7950 800 7966 856
rect 8318 800 8334 856
rect 8686 800 8702 856
rect 9054 800 9070 856
rect 9422 800 9438 856
rect 9790 800 9806 856
rect 10158 800 10174 856
rect 10526 800 10542 856
rect 10894 800 10910 856
rect 11354 800 11370 856
rect 11722 800 11738 856
rect 12090 800 12106 856
rect 12458 800 12474 856
rect 12826 800 12842 856
rect 13194 800 13210 856
rect 13562 800 13578 856
rect 13930 800 13946 856
rect 14298 800 14314 856
rect 14666 800 14682 856
rect 15126 800 15142 856
rect 15494 800 15510 856
rect 15862 800 15878 856
rect 16230 800 16246 856
rect 16598 800 16614 856
rect 16966 800 16982 856
rect 17334 800 17350 856
rect 17702 800 17718 856
rect 18070 800 18086 856
rect 18438 800 18454 856
rect 18898 800 18914 856
rect 19266 800 19282 856
rect 19634 800 19650 856
rect 20002 800 20018 856
rect 20370 800 20386 856
rect 20738 800 20754 856
rect 21106 800 21122 856
rect 21474 800 21490 856
rect 21842 800 21858 856
rect 22210 800 22226 856
rect 22670 800 22686 856
rect 23038 800 23054 856
rect 23406 800 23422 856
rect 23774 800 23790 856
rect 24142 800 24158 856
rect 24510 800 24526 856
rect 24878 800 24894 856
rect 25246 800 25262 856
rect 25614 800 25630 856
rect 25982 800 25998 856
rect 26442 800 26458 856
rect 26810 800 26826 856
rect 27178 800 27194 856
rect 27546 800 27562 856
rect 27914 800 27930 856
rect 28282 800 28298 856
rect 28650 800 28666 856
rect 29018 800 29034 856
rect 29386 800 29402 856
rect 29754 800 29770 856
rect 30214 800 30230 856
rect 30582 800 30598 856
rect 30950 800 30966 856
rect 31318 800 31334 856
rect 31686 800 31702 856
rect 32054 800 32070 856
rect 32422 800 32438 856
rect 32790 800 32806 856
rect 33158 800 33174 856
rect 33526 800 33542 856
rect 33986 800 34002 856
rect 34354 800 34370 856
rect 34722 800 34738 856
rect 35090 800 35106 856
rect 35458 800 35474 856
rect 35826 800 35842 856
rect 36194 800 36210 856
rect 36562 800 36578 856
rect 36930 800 36946 856
rect 37298 800 37314 856
rect 37758 800 37774 856
rect 38126 800 38142 856
rect 38494 800 38510 856
rect 38862 800 38878 856
rect 39230 800 39246 856
rect 39598 800 39614 856
rect 39966 800 39982 856
rect 40334 800 40350 856
rect 40702 800 40718 856
rect 41070 800 41086 856
rect 41530 800 41546 856
rect 41898 800 41914 856
rect 42266 800 42282 856
rect 42634 800 42650 856
rect 43002 800 43018 856
rect 43370 800 43386 856
rect 43738 800 43754 856
rect 44106 800 44122 856
rect 44474 800 44490 856
rect 44842 800 44858 856
rect 45302 800 45318 856
rect 45670 800 45686 856
rect 46038 800 46054 856
rect 46406 800 46422 856
rect 46774 800 46790 856
rect 47142 800 47158 856
rect 47510 800 47526 856
rect 47878 800 47894 856
rect 48246 800 48262 856
rect 48614 800 48630 856
rect 49074 800 49090 856
rect 49442 800 49458 856
rect 49810 800 49826 856
rect 50178 800 50194 856
rect 50546 800 50562 856
rect 50914 800 50930 856
rect 51282 800 51298 856
rect 51650 800 51666 856
rect 52018 800 52034 856
rect 52386 800 52402 856
rect 52846 800 52862 856
rect 53214 800 53230 856
rect 53582 800 53598 856
rect 53950 800 53966 856
rect 54318 800 54334 856
rect 54686 800 54702 856
rect 55054 800 55070 856
rect 55422 800 55438 856
rect 55790 800 55806 856
rect 56158 800 56174 856
rect 56618 800 56634 856
rect 56986 800 57002 856
rect 57354 800 57370 856
rect 57722 800 57738 856
rect 58090 800 58106 856
rect 58458 800 58474 856
rect 58826 800 58842 856
rect 59194 800 59210 856
rect 59562 800 59578 856
<< obsm3 >>
rect 3049 2143 57119 38997
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
<< obsm4 >>
rect 9811 37664 33797 38997
rect 9811 26963 19488 37664
rect 19968 26963 33797 37664
<< labels >>
rlabel metal2 s 202 39200 258 40000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 15934 39200 15990 40000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 17498 39200 17554 40000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 19062 39200 19118 40000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 20718 39200 20774 40000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 22282 39200 22338 40000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 23846 39200 23902 40000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25410 39200 25466 40000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 26974 39200 27030 40000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28538 39200 28594 40000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30194 39200 30250 40000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 1766 39200 1822 40000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31758 39200 31814 40000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 33322 39200 33378 40000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34886 39200 34942 40000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 36450 39200 36506 40000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 38014 39200 38070 40000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 39578 39200 39634 40000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 41234 39200 41290 40000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 42798 39200 42854 40000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 44362 39200 44418 40000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45926 39200 45982 40000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3330 39200 3386 40000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 47490 39200 47546 40000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 49054 39200 49110 40000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 50710 39200 50766 40000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 52274 39200 52330 40000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53838 39200 53894 40000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 55402 39200 55458 40000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 56966 39200 57022 40000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 58530 39200 58586 40000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 4894 39200 4950 40000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6458 39200 6514 40000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 8022 39200 8078 40000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 9586 39200 9642 40000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 11242 39200 11298 40000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 12806 39200 12862 40000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 14370 39200 14426 40000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 662 39200 718 40000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 16486 39200 16542 40000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 18050 39200 18106 40000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 19614 39200 19670 40000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 21178 39200 21234 40000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 22742 39200 22798 40000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 24398 39200 24454 40000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 25962 39200 26018 40000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 27526 39200 27582 40000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29090 39200 29146 40000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30654 39200 30710 40000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 2226 39200 2282 40000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32218 39200 32274 40000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33874 39200 33930 40000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 35438 39200 35494 40000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 37002 39200 37058 40000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 38566 39200 38622 40000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 40130 39200 40186 40000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 41694 39200 41750 40000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 43258 39200 43314 40000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 44914 39200 44970 40000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 46478 39200 46534 40000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 3882 39200 3938 40000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 48042 39200 48098 40000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 49606 39200 49662 40000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 51170 39200 51226 40000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 52734 39200 52790 40000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 54390 39200 54446 40000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 55954 39200 56010 40000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 57518 39200 57574 40000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 59082 39200 59138 40000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5446 39200 5502 40000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 7010 39200 7066 40000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 8574 39200 8630 40000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 10138 39200 10194 40000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 11702 39200 11758 40000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 13266 39200 13322 40000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 14922 39200 14978 40000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1214 39200 1270 40000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 17038 39200 17094 40000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 18602 39200 18658 40000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 20166 39200 20222 40000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 21730 39200 21786 40000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23294 39200 23350 40000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 24858 39200 24914 40000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 26422 39200 26478 40000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28078 39200 28134 40000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 29642 39200 29698 40000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31206 39200 31262 40000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 2778 39200 2834 40000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32770 39200 32826 40000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 34334 39200 34390 40000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35898 39200 35954 40000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 37554 39200 37610 40000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 39118 39200 39174 40000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 40682 39200 40738 40000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42246 39200 42302 40000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 43810 39200 43866 40000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 45374 39200 45430 40000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 47030 39200 47086 40000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4342 39200 4398 40000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 48594 39200 48650 40000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50158 39200 50214 40000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 51722 39200 51778 40000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 53286 39200 53342 40000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 54850 39200 54906 40000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56414 39200 56470 40000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 58070 39200 58126 40000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 59634 39200 59690 40000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 5906 39200 5962 40000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 7562 39200 7618 40000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 9126 39200 9182 40000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 10690 39200 10746 40000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 12254 39200 12310 40000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 13818 39200 13874 40000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15382 39200 15438 40000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 503 nsew ground input
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 662 0 718 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 40000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 2759564
string GDS_START 267730
<< end >>

